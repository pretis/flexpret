module Top(
  output [7:0] LEDS
);

  assign LEDS = 8'b01010101;
  
endmodule
